library verilog;
use verilog.vl_types.all;
entity MIPSTestBench is
end MIPSTestBench;
